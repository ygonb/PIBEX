CircuitMaker Text
5.6
Probes: 3
S1_1
AC Analysis
0 709 257 65280
S1_1
Transient Analysis
0 711 257 65280
S1_2
Transient Analysis
1 429 257 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 140 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1532 489
9961490 0
0
6 Title:
5 Name:
0
0
0
12
12 SPDT Switch~
164 679 257 0 3 11
0 3 5 3
0
0 0 4720 0
0
2 S1
-7 -15 7 -7
0
0
0
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
0 0 0 0 1 0 0 0
1 S
9197 0 0
2
43916.7 0
0
7 Ground~
168 321 330 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9624 0 0
2
43916.7 1
0
11 Signal Gen~
195 276 309 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1176256512 0 1036831949
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 18
20
1 10000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -100m/100mV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(0 100m 10k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3383 0 0
2
43916.7 2
0
7 summer~
219 379 256 0 3 7
0 7 6 5
0
0 0 50000 0
3 SUM
-4 -31 17 -23
2 U2
0 -41 14 -33
0
0
16 %D [%1 %2] %3 %M
0
11 type:summer
0
7

0 0 0 0 0 0 0 0
65 0 0 0 1 0 0 0
1 U
8868 0 0
2
43916.7 3
0
11 Signal Gen~
195 272 222 0 64 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1114636288 1075838976 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 60 2.5 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 1.5/3.5V
-28 -30 28 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(2.5 1 60 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3645 0 0
2
43916.7 4
0
7 Ground~
168 317 243 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8552 0 0
2
43916.7 5
0
10 Op-Amp5:A~
219 567 264 0 5 11
0 8 3 10 11 3
0
0 0 848 0
5 LM324
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 512 1 0 0 0
1 U
3924 0 0
2
43916.7 6
0
10 Capacitor~
219 513 312 0 2 5
0 3 9
0
0 0 848 180
5 .47uF
-17 -18 18 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8841 0 0
2
43916.7 7
0
7 Ground~
168 562 188 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4326 0 0
2
43916.7 8
0
10 Capacitor~
219 539 223 0 2 5
0 8 2
0
0 0 848 90
5 .47uF
5 0 40 8
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4303 0 0
2
43916.7 9
0
9 Resistor~
219 453 256 0 2 5
0 5 9
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
651 0 0
2
43916.7 10
0
9 Resistor~
219 508 256 0 2 5
0 9 8
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5592 0 0
2
43916.7 11
0
15
1 0 3 0 0 4224 0 1 0 0 0 2
696 257
725 257
3 0 3 0 0 8192 4 1 0 0 11 3
662 261
662 264
624 264
0 2 5 0 0 8320 0 0 1 6 0 5
427 256
427 154
650 154
650 253
662 253
1 2 6 0 0 8320 0 3 4 0 0 4
307 304
341 304
341 265
355 265
2 1 2 0 0 4096 0 3 2 0 0 3
307 314
321 314
321 324
3 1 5 0 0 0 0 4 11 0 0 2
417 256
435 256
1 1 7 0 0 4224 0 5 4 0 0 4
303 217
342 217
342 247
355 247
2 1 2 0 0 0 0 5 6 0 0 3
303 227
317 227
317 237
2 1 2 0 0 4224 0 10 9 0 0 4
539 214
539 169
562 169
562 182
1 0 8 0 0 4224 0 10 0 0 14 2
539 232
539 256
0 5 3 0 0 4224 4 0 7 12 0 4
540 312
624 312
624 264
585 264
2 1 3 0 0 0 4 7 8 0 0 4
549 270
540 270
540 312
522 312
2 0 9 0 0 8320 0 8 0 0 15 3
504 312
482 312
482 256
2 1 8 0 0 0 0 12 7 0 0 4
526 256
541 256
541 258
549 258
2 1 9 0 0 0 0 11 12 0 0 2
471 256
490 256
0
0
25 0 1
0
0
0
0 0 0
0
0 0 0
1000 1 1 10000
0 0.05 5e-07 5e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
